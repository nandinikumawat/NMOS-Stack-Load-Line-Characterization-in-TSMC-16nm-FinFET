** Generated for: hspiceD
** Generated on: Oct 27 21:09:02 2025
** Design library name: ee8310
** Design cell name: NMOS_stack
** Design view name: schematic

** Library name: ee8310
** Cell name: NMOS_stack
** View name: schematic
xm1 vx b vss vss nch_svt_mac l=16e-9 nfin=2 w=58e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm0 vdd a vx vss nch_svt_mac l=16e-9 nfin=2 w=58e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
.END

